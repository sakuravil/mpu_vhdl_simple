library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity clkgen is
end clkgen;

architecture Behavioral of clkgen is

begin


end Behavioral;

